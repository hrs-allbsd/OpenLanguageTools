Ang.
Ank.
Avd.
Avg.
Avs.
Betr.
Bil.
Bitr.
Bull.
Dir.
Dvs.
Enl.
Exp.
Exv.
F�lj.
Fr.
Fr.o.m.
F�reg.
Gm.
Hr.
Kl.
Mag.
Prof.
T.ex.
Tel.
U.S.
U.S.A.
ang.
ank.
avd.
avg.
avs.
betr.
bil.
bitr.
bull.
dir.
dr.
dvs.
enl.
exp.
exv.
f�lj.
fr.
fr.o.m.
f�reg.
gm.
hr.
kl.
mag.
prof.
t.ex.
tel.
Adr.
adr.
Bl.a.
bl.a.
Civ.ek.
civ.ek.
Civ.ing.
civ.ing.
Co.
Div.
div.
Doc.
doc.
E.dyl.
e.dyl.
el.
etc.
Ev.
ev.
Ex.
ex.
Exkl.
exkl.
F.d.
f.d.
ff.
Forts.
forts.
F.�.
f.�.
Ibl.
ibl.
Inkl.
inkl.
I st.f.
i st.f.
Kr.
kr.
lev.
Max.
max.
M.fl.
m.fl.
Min.
min.
m.m.
Nuv.
nuv.
Obs.
obs.
o.d.
o.dyl.
Ordf.
ordf.
osv.
Pg.
pg.
pl.
plur.
P.S.
Sek.
sek.
Sekr.
sekr.
Sid.
sid.
Sign.
sign.
s.k.
Spec.
spec.
St.
st.
tekn.
Tf.
tf.
Tim.
tim.
tr.
T.v.
t.v.
Ung.
ung.
Uppl.
uppl.
v.
Vol.
vol.
�rg.
�rg.
�v.
�.
